** sch_path: /foss/designs/ihp-inverter/xschem/tb_inverter.sch
**.subckt tb_inverter
VIN vin GND PULSE(0 3 0 1n 1n 4n 10n)
VDD vdd GND 3
x1 vdd vin vout_sim GND inverter
x2 vdd vin vout_kl GND inverter_ext
**** begin user architecture code

.lib cornerMOShv.lib mos_tt





.include tb_inverter.save
.param temp=27
.control
save all
op
tran 10p 20n
write tb_inverter.raw
.endc



.inc /foss/designs/ihp-inverter/klayout/inverter_ext.spice

**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /foss/designs/ihp-inverter/xschem/inverter.sym
** sch_path: /foss/designs/ihp-inverter/xschem/inverter.sch
.subckt inverter VDD A Y VSS
*.ipin A
*.opin Y
*.iopin VDD
*.iopin VSS
XM1 Y A VSS VSS sg13_hv_nmos w=0.3u l=0.45u ng=1 m=1
XM2 Y A VDD VDD sg13_hv_pmos w=0.3u l=0.45u ng=1 m=1
.ends

.GLOBAL GND
.end
